module and_gate (a,b,c);
//  declaring inputs and output
 input a;
 input b;

 output c;

// defining bits to  input [31:0] D;
 
//  Gate level modeling
 
 and a1 (c,a,b);


endmodule
